//=============================================================================
// File: pkt_proc_scoreboard_new.sv
// Description: New Simple Packet Processor UVM Scoreboard
// Author: Assistant
// Date: 2024
//=============================================================================


class pkt_proc_scoreboard extends uvm_scoreboard;
    `uvm_component_utils(pkt_proc_scoreboard)

    uvm_analysis_imp #(pkt_proc_seq_item, pkt_proc_scoreboard) analysis_export;

    // Configuration parameters (matching RTL)
    parameter int DEPTH = 16384;
    parameter int PCK_LEN_DEPTH = 32;
    parameter int DATA_WIDTH = 32;
    parameter int ADDR_WIDTH = 14;
    parameter int PCK_LEN = 12;

    // Reference model state machines (matching RTL)
    typedef enum {IDLE_W, WRITE_HEADER, WRITE_DATA} write_state_e;
    typedef enum {IDLE_R, READ_HEADER, READ_DATA} read_state_e;
    
    write_state_e write_state;
    write_state_e write_state_next; // next-state mirror for write FSM
    read_state_e read_state;
    read_state_e read_state_next; // mirror RTL present/next state split
    read_state_e read_state_prev; // previous state for output generation timing
    
    // Reference model internal state
    bit [31:0] ref_buffer[0:16383];  // Main buffer
    bit [11:0] ref_pck_len_buffer[0:31];  // Packet length buffer
    // Buffer state tracking
    bit [14:0] ref_wr_ptr;           // Write pointer (address) - CRITICAL for concurrent operations
    bit [14:0] ref_wr_ptr_next;      // Next write pointer
    bit [14:0] ref_rd_ptr;           // Read pointer (for buffer reads)
    bit [11:0] ref_pck_len_wr_ptr;   // Packet length FIFO write pointer
    bit [11:0] ref_pck_len_rd_ptr;   // Packet length FIFO read pointer
    bit [14:0] ref_wr_lvl;           // Write level (matching RTL output)
    bit [11:0] ref_count_r;          // Read counter (matching RTL count_r)
    
    // Packet length tracking
    bit [11:0] ref_packet_length;      // Current packet length (from read path)
    bit [11:0] ref_packet_length_w;    // Write path packet length (for pck_invalid checks)
    bit [11:0] ref_count_w_prev;       // Previous cycle's count_w for packet drop calculations
    bit [11:0] ref_count_w2_prev;      // Previous cycle's count_w2 for packet drop calculations
    bit [11:0] ref_count_w;            // Current cycle's count_w value
    bit [11:0] ref_count_w_next;       // Next cycle's count_w value (for proper timing)
    bit [11:0] ref_count_w2;           // Second count_w variable (matching new RTL)
    bit [11:0] ref_count_w2_next;      // Next cycle's count_w2 value
    bit ref_buffer_full, ref_buffer_empty;
    bit ref_pck_len_full, ref_pck_len_empty;
    bit ref_pck_proc_overflow, ref_pck_proc_underflow;
    bit ref_packet_drop;
    bit ref_packet_drop_prev;  // track rising edge of packet_drop for debug
    bit invalid_1, invalid_3, invalid_4, invalid_5, invalid_6, any_invalid_condition; // packet drop conditions
    
    // Expected outputs
    bit ref_out_sop, ref_out_eop;
    bit [31:0] ref_rd_data_o;
    bit ref_pck_proc_almost_full, ref_pck_proc_almost_empty;
    
    // Pipeline registers (matching RTL exactly)
    bit ref_in_sop_r, ref_in_sop_r1, ref_in_sop_r2;
    bit ref_in_eop_r, ref_in_eop_r1, ref_in_eop_r2;
    bit ref_enq_req_r, ref_enq_req_r1;
    bit [31:0] ref_wr_data_r, ref_wr_data_r1;
    bit ref_pck_len_valid_r, ref_pck_len_valid_r1;
    bit [11:0] ref_pck_len_i_r, ref_pck_len_i_r1;
    bit ref_deq_req_r;   // registered deq_req (1-cycle delayed)
    bit ref_deq_req_r1;  // sampling stage for deq_req
    
    // Additional signals
    bit ref_empty_de_assert;
    bit ref_buffer_empty_r;
    bit ref_wr_en, ref_rd_en;
    bit ref_wr_en_prev;  // Previous cycle's write enable
    bit ref_rd_en_prev;  // Previous cycle's read enable
    bit ref_deq_req_prev;  // Previous cycle's dequeue request (for out_sop timing)
    
    // Read pipeline delay (matching DUT timing)
    //bit [31:0] ref_rd_data_delayed;  // Delayed read data output
    bit ref_deq_req_prev2;  // Two cycles ago dequeue request (for out_sop timing)
    bit ref_buffer_full_prev;   // Previous cycle's buffer_full
    bit ref_buffer_empty_prev;  // Previous cycle's buffer_empty
    
    // CRITICAL FIX: Add two-cycle delayed buffer_full for overflow detection
    // Overflow should go high AFTER one clock pulse after pck_proc_full goes high
    bit ref_buffer_full_prev2;  // Two cycles ago buffer_full (for overflow timing)
    
    // CRITICAL FIX: Add read pointer next value for proper timing alignment
    bit [13:0] ref_rd_ptr_next;  // Next cycle's read pointer (for 1-cycle delay matching DUT)
    
    // Write level tracking (matching RTL's always_ff behavior)
    bit [14:0] ref_wr_lvl_next;     // Next cycle's wr_lvl value (15 bits: [ADDR_WIDTH:0])
    bit ref_overflow;               // Internal overflow signal (matching int_buffer_top)
    bit ref_overflow_prev;          // Previous cycle's overflow
    bit ref_reset_active;           // Flag to track if reset is currently active
    
    // One-cycle delayed signals (matching RTL's always_ff outputs)
    bit ref_buffer_empty_delayed;   // One-cycle delayed buffer_empty
    
    // Temporary variables for combinational calculations
    bit temp_full, temp_empty;
    
    // Statistics
    int total_transactions = 0;
    int errors = 0;

    bit data_available;
    bit data_available_next;
    bit data_available_for_comparison;



    function new(string name, uvm_component parent);
        super.new(name, parent);
        analysis_export = new("analysis_export", this);
        initialize_reference_model();
    endfunction

    function void initialize_reference_model();
        // Initialize state machines
        write_state = IDLE_W;
        write_state_next = IDLE_W;
        read_state = IDLE_R;
        read_state_next = IDLE_R;
        read_state_prev = IDLE_R;  // Initialize previous state
        
        // Initialize pointers and counters
        ref_wr_ptr = 0;           // Write pointer starts at 0
        ref_wr_ptr_next = 0;      // Next write pointer starts at 0
        ref_rd_ptr = 0;
        ref_rd_ptr_next = 0;  // Initialize next cycle's read pointer
        ref_pck_len_wr_ptr = 0;
        ref_pck_len_rd_ptr = 0;
        ref_wr_lvl = 0;
        ref_count_w = 0;            // Current count_w starts at 0
        ref_count_w_next = 0;       // Next count_w starts at 0
        ref_count_w_prev = 0;       // Initialize previous count_w
        ref_count_w2 = 0;           // Second count_w starts at 0
        ref_count_w2_next = 0;      // Next count_w2 starts at 0
        ref_count_w2_prev = 0;      // Initialize previous count_w2
        ref_count_r = 0;
        ref_packet_length = 0;
        ref_packet_length_w = 0;
        `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: ref_packet_length_w initialized to 0", $time), UVM_LOW)
        
        // Initialize buffer states
        ref_buffer_full = 0;
        ref_buffer_empty = 1;
        ref_pck_len_full = 0;
        ref_pck_len_empty = 1;
        

        // Initialize flags
        ref_pck_proc_overflow = 0;
        ref_pck_proc_underflow = 0;
        ref_packet_drop = 0;
        ref_packet_drop_prev = 0;
        invalid_1 = 0;
        invalid_3 = 0;
        invalid_4 = 0;
        invalid_5 = 0;
        invalid_6 = 0;
        any_invalid_condition = 0;
        
        // Initialize outputs
        ref_out_sop = 0;
        ref_out_eop = 0;
        ref_rd_data_o = 0;
        ref_pck_proc_almost_full = 0;
        ref_pck_proc_almost_empty = 0;
        
        // Initialize pipeline registers
        ref_in_sop_r = 0; ref_in_sop_r1 = 0; ref_in_sop_r2 = 0;
        ref_in_eop_r = 0; ref_in_eop_r1 = 0; ref_in_eop_r2 = 0;
        ref_enq_req_r = 0; ref_enq_req_r1 = 0;
        ref_wr_data_r = 0; ref_wr_data_r1 = 0;
        ref_pck_len_valid_r = 0; ref_pck_len_valid_r1 = 0;
        ref_pck_len_i_r = 0; ref_pck_len_i_r1 = 0;
        ref_deq_req_r = 0;
        
        // Initialize additional signals
        ref_empty_de_assert = 1;
        ref_buffer_empty_r = 1;
        ref_wr_en = 0;
        ref_rd_en = 0;
        ref_wr_en_prev = 0;
        ref_rd_en_prev = 0;
        ref_deq_req_prev = 0;
        //ref_rd_data_delayed = 0;
        ref_deq_req_prev2 = 0;
        ref_buffer_full_prev = 0;
        ref_buffer_empty_prev = 1;
        ref_buffer_full_prev2 = 0;  // Initialize two-cycle delayed buffer_full
        
        // Initialize write level tracking
        ref_wr_lvl_next = 0;
        ref_overflow = 0;
        ref_overflow_prev = 0;
        
        // Initialize delayed signals
        ref_buffer_empty_delayed = 1;
        
        // Initialize reset flag
        ref_reset_active = 0;
        
        // Initialize temporary variables
        temp_full = 0;
        temp_empty = 0;

        data_available = 0;
        data_available_next = 0;
        data_available_for_comparison = 0;
    endfunction

    function void write(pkt_proc_seq_item tr);
        total_transactions++;
        
        `uvm_info("SCOREBOARD_NEW", $sformatf("Processing transaction #%0d", total_transactions), UVM_LOW)
        
        // All transactions are now clock-based - unified processing
        `uvm_info("CLOCK_EDGE_TRANSACTION", $sformatf("Time=%0t: Processing clock edge transaction", $time), UVM_LOW)
        
        // Update reference model (includes packet drop detection and all other logic)
        update_reference_model(tr);
        
        // Compare outputs with DUT
        compare_outputs(tr);
        
        // Update wr_lvl and count_w for next cycle (matching RTL always_ff timing)
        if (ref_wr_lvl_next != ref_wr_lvl) begin
            `uvm_info("WR_LVL_UPDATE", $sformatf("Time=%0t: Updating wr_lvl after comparison: %0d -> %0d (for next cycle)", 
                     $time, ref_wr_lvl, ref_wr_lvl_next), UVM_LOW)
            ref_wr_lvl = ref_wr_lvl_next;
        end
        if (ref_count_w_next != ref_count_w) begin
            `uvm_info("COUNT_W_UPDATE", $sformatf("Time=%0t: Updating count_w after comparison: %0d -> %0d (for next cycle)", 
                     $time, ref_count_w, ref_count_w_next), UVM_LOW)
            ref_count_w = ref_count_w_next;
        end
        
        // CRITICAL FIX: Update count_w2 to match new RTL implementation
        if (ref_count_w2_next != ref_count_w2) begin
            `uvm_info("COUNT_W2_UPDATE", $sformatf("Time=%0t: Updating count_w2 after comparison: %0d -> %0d (for next cycle)", 
                     $time, ref_count_w2, ref_count_w2_next), UVM_LOW)
            ref_count_w2 = ref_count_w2_next;
        end
    endfunction

    function void update_reference_model(pkt_proc_seq_item tr);
        // ============================================================================
        // CORRECT EXECUTION ORDER - Resolving ALL Dependencies
        // ============================================================================
        // 
        // RTL Reality:
        // - ALL always_ff blocks execute simultaneously at posedge clock using <=
        // - Combinational logic (always_comb) executes continuously
        // - State updates happen at clock edge using values from previous cycle
        //
        // Scoreboard Emulation:
        // - Use CURRENT pipeline register values for current cycle logic (matching RTL)
        // - Update all state variables simultaneously at end (matching RTL <= behavior)
        // - Ensure combinational logic uses consistent values from same cycle
        //
        // Key Principle: Each function uses values that would be available in RTL
        // at the start of the clock cycle, not values calculated during the cycle
        // ============================================================================
        
        // Debug current states being processed
        `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: Processing with states - WRITE: %0d, READ: %0d", 
                 $time, write_state, read_state), UVM_LOW)
        
        // ============================================================================
        // PHASE 1: Reset logic (highest priority)
        // ============================================================================
        handle_reset_logic(tr);                    // Sets ref_reset_active
        
        // ref_buffer_full_prev2 = ref_buffer_full_prev;  // Two-cycle delay for overflow
        // ref_buffer_full_prev  = ref_buffer_full;
        // ref_buffer_empty_prev = ref_buffer_empty;
        // ref_overflow_prev = ref_overflow;

        // ============================================================================
        // PHASE 16: Buffer synchronization
        // ============================================================================
        // CRITICAL FIX: Calculate wr_lvl_next based on NEXT cycle's pointers (matching RTL exactly)
        // RTL: wr_lvl = wr_ptr - rd_ptr, but pointers update with 1-cycle delay
        // So for current cycle: wr_lvl_next = wr_ptr_next - rd_ptr_next

        // ref_wr_lvl_next = ref_wr_ptr_next - ref_rd_ptr_next;
        // `uvm_info("WR_LVL_NEXT", $sformatf("Time=%0t: wr_lvl_next=%0d, wr_ptr_next=%0d, rd_ptr_next=%0d", $time, ref_wr_lvl_next, ref_wr_ptr_next, ref_rd_ptr_next), UVM_LOW)
        // CRITICAL FIX: Update pointers for next cycle (matching RTL always_ff behavior)
        ref_wr_ptr = ref_wr_ptr_next;  // Update write pointer
        ref_rd_ptr = ref_rd_ptr_next;  // Update read pointer
        
        // CRITICAL FIX: Update wr_lvl for next cycle (matching RTL always_ff behavior)
        ref_wr_lvl = ref_wr_lvl_next;

        ref_buffer_full_prev  = ref_buffer_full;
        ref_buffer_empty_prev = ref_buffer_empty;
        ref_overflow_prev = ref_overflow;
        ref_buffer_full_prev2 = ref_buffer_full_prev;  // Two-cycle delay for overflow
        
        // ============================================================================
        // PHASE 2: Update buffer states FIRST (before packet drop logic)
        // ============================================================================
        update_buffer_states();                    // Sets ref_buffer_full, ref_buffer_empty
        
        // Debug current cycle inputs for state transitions
        `uvm_info("STATE_INPUTS", $sformatf("Time=%0t: Current inputs - in_sop=%0b, in_eop=%0b, enq_req=%0b, pck_len_valid=%0b, pck_len_i=%0d", 
                 $time, tr.in_sop, tr.in_eop, tr.enq_req, tr.pck_len_valid, tr.pck_len_i), UVM_LOW)
        
        // ============================================================================
        // PHASE 3: Update combinational outputs (uses updated buffer states)
        // ============================================================================
        update_combinational_outputs(tr);          // Sets ref_pck_proc_* outputs
        
        // ============================================================================
        // PHASE 4: Update internal overflow (uses updated buffer states)
        // ============================================================================
        update_internal_overflow();                // Sets ref_overflow
        
        // ============================================================================
        // PHASE 5: Update packet drop logic FIRST (before enable generation)
        // ============================================================================
        update_packet_drop_logic(tr);              // Sets ref_packet_drop
        
        // Handle packet drop logic for count_w_next
        if (ref_packet_drop) begin
            `uvm_info("PKT_DROP_DEBUG", $sformatf("Time=%0t: PACKET_DROP detected: count_w=%0d, wr_lvl=%0d", 
                     $time, ref_count_w, ref_wr_lvl), UVM_LOW)
            
            // CRITICAL FIX: RTL uses always_ff, so wr_lvl updates at NEXT clock edge
            // The wr_lvl_next calculation is handled in update_write_level_next()
            // Here we just calculate count_w_next for next packet (matching RTL)
            ref_count_w_next = 0;
            
            `uvm_info("PKT_DROP_DEBUG", $sformatf("Time=%0t: PACKET_DROP: count_w_next set to 0, wr_lvl_next will be calculated in update_write_level_next()", 
                     $time), UVM_LOW)
        end
        
        // CRITICAL FIX: Add count_w2 logic to match new RTL implementation
        // New RTL has different reset logic for count_w2
        if (ref_packet_drop) begin
            if (ref_in_sop_r1 && !ref_in_eop_r1) begin
                // Special case: in_sop_r1 && !in_eop_r1 && packet_drop
                ref_count_w2_next = 1;
                `uvm_info("COUNT_W2_DEBUG", $sformatf("Time=%0t: COUNT_W2 special case: in_sop_r1=%0b, in_eop_r1=%0b, packet_drop=%0b, count_w2_next=1", 
                         $time, ref_in_sop_r1, ref_in_eop_r1, ref_packet_drop), UVM_LOW)
            end else begin
                // Normal packet drop: reset count_w2 to 0
                ref_count_w2_next = 0;
                `uvm_info("COUNT_W2_DEBUG", $sformatf("Time=%0t: COUNT_W2 normal reset: count_w2_next=0", $time), UVM_LOW)
            end
        end else if (ref_in_eop_r1 && (write_state == WRITE_DATA)) begin
            // Packet completed normally: reset count_w2 to 0
            ref_count_w2_next = 0;
            `uvm_info("COUNT_W2_DEBUG", $sformatf("Time=%0t: COUNT_W2 packet complete: count_w2_next=0", $time), UVM_LOW)
        end else if (ref_wr_en && !ref_buffer_full) begin
            // Successful write: increment count_w2
            ref_count_w2_next = ref_count_w2 + 1;
            `uvm_info("COUNT_W2_DEBUG", $sformatf("Time=%0t: COUNT_W2 increment: count_w2=%0d -> %0d", 
                     $time, ref_count_w2, ref_count_w2_next), UVM_LOW)
        end else begin
            // No change
            ref_count_w2_next = ref_count_w2;
        end
        
        // ============================================================================
        // PHASE 6: Generate enables (uses packet drop and current states)
        // ============================================================================
        generate_write_read_enables(tr);           // Uses ref_packet_drop, sets ref_wr_en, ref_rd_en
         
        // ref_buffer_full_prev  = ref_buffer_full;
        // //ref_buffer_empty_prev = ref_buffer_empty;
        // ref_overflow_prev = ref_overflow;
        // ref_buffer_full_prev2 = ref_buffer_full_prev;  // Two-cycle delay for overflow
        
       
        // ============================================================================
        // PHASE 7: Update write level (uses packet drop, buffer states, and enables)
        // ============================================================================
        update_write_level_next();                 // Uses ref_packet_drop, ref_buffer_full, ref_buffer_empty
        
        // CRITICAL FIX: Update buffer states AFTER buffer operations (matching RTL timing)
        // This ensures ref_buffer_empty reflects the current state after reads/writes
        update_combinational_outputs(tr);
        
        // ============================================================================
        // PHASE 8: Buffer operations (uses correct enables, write level, and packet drop)
        // ============================================================================
        if (!ref_packet_drop) begin
            // Write operations - only when packet is valid
            if (ref_wr_en && !ref_buffer_full) begin
                // CRITICAL DEBUG: Track buffer writes when wr_lvl = 0
                if (ref_wr_lvl == 0) begin
                    `uvm_info("BUFFER_WRITE_DEBUG", $sformatf("Time=%0t: WRITING TO BUFFER[0]: wr_en=%0b, buffer_full=%0b, state=%0d, data=0x%0h", 
                             $time, ref_wr_en, ref_buffer_full, write_state, ref_wr_data_r), UVM_LOW)
                end
                
                if (write_state == WRITE_HEADER) begin
                    ref_buffer[ref_wr_ptr[13:0]] = ref_wr_data_r;  // Use write pointer, NOT wr_lvl
                end else if (write_state == WRITE_DATA) begin
                    ref_buffer[ref_wr_ptr[13:0]] = ref_wr_data_r;  // Use write pointer, NOT wr_lvl
                end
                
                // CRITICAL FIX: Increment write pointer for successful write operations
                ref_wr_ptr_next = ref_wr_ptr + 1;
                
                // CRITICAL FIX: Increment count_w_next for successful write operations
                ref_count_w_next = ref_count_w + 1;
                `uvm_info("COUNT_W_DEBUG", $sformatf("Time=%0t: count_w_next set to %0d (state=%0d, wr_en=%0b, wr_ptr=%0d->%0d, buffer[%0d]=0x%0h)", 
                         $time, ref_count_w_next, write_state, ref_wr_en, ref_wr_ptr, ref_wr_ptr_next, ref_wr_ptr[13:0], ref_wr_data_r1), UVM_LOW)
            end
            
            // CRITICAL FIX: Packet length buffer operations (matching RTL exactly)
            // RTL writes to pck_len_buffer in WRITE_HEADER state regardless of wr_en
            if (write_state == WRITE_HEADER) begin
                // Use RTL logic exactly: pck_len_r2 = (pck_len_valid_r1) ? pck_len_i_r1 : ((in_sop_r1) ? wr_data_r1[11:0] : packet_length)
                // CRITICAL: These _r1 values contain the PREVIOUS cycle's values (when in_sop=1, pck_len_valid=1)
                bit [11:0] pck_len_r2_value;
                if (ref_pck_len_valid_r1) begin
                    pck_len_r2_value = ref_pck_len_i_r1;
                    `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: WRITE_HEADER: Using pck_len_i_r1=%0d (pck_len_valid_r1=1)", 
                             $time, ref_pck_len_i_r1), UVM_LOW)
                end else if (ref_in_sop_r1) begin
                    pck_len_r2_value = ref_wr_data_r1[11:0];
                    `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: WRITE_HEADER: Using wr_data_r1[11:0]=%0d (in_sop_r1=1)", 
                             $time, ref_wr_data_r1[11:0]), UVM_LOW)
                end else begin
                    pck_len_r2_value = ref_packet_length_w;  // Keep previous value
                    `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: WRITE_HEADER: Using prev_packet_length=%0d (both conditions false)", 
                             $time, ref_packet_length_w), UVM_LOW)
                end
                
                // Write to packet length buffer (matching RTL pck_len_wr_en = 1'b1 in WRITE_HEADER)
                ref_pck_len_buffer[ref_pck_len_wr_ptr[4:0]] = pck_len_r2_value;
                ref_pck_len_wr_ptr = ref_pck_len_wr_ptr + 1;
                
                // Update write-path packet length mirror for pck_invalid checks
                ref_packet_length_w = pck_len_r2_value;
                
                // Debug print for packet length assignment
                `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: WRITE_HEADER: pck_len_r2=%0d (pck_len_valid_r1=%0b, in_sop_r1=%0b, pck_len_i_r1=%0d, wr_data_r1[11:0]=%0d, prev_packet_length=%0d)", 
                         $time, pck_len_r2_value, ref_pck_len_valid_r1, ref_in_sop_r1, ref_pck_len_i_r1, ref_wr_data_r1[11:0], ref_packet_length_w), UVM_LOW)
            end
        end else begin
            // CRITICAL FIX: When packet drop is detected, adjust write pointer (matching RTL exactly)
            // RTL: wr_ptr <= wr_ptr - count_w (or wr_ptr - count_w + 1 for invalid_3)
            if (invalid_3) begin
                // Special case: pck_drop && invalid_3
                ref_wr_ptr_next = ref_wr_ptr - ref_count_w + 1;
                `uvm_info("PKT_DROP_DEBUG", $sformatf("Time=%0t: Packet drop (invalid_3): wr_ptr %0d -> %0d (count_w=%0d, +1)", 
                         $time, ref_wr_ptr, ref_wr_ptr_next, ref_count_w), UVM_LOW)
            end else begin
                // Normal packet drop: decrement wr_ptr by count_w
                ref_wr_ptr_next = ref_wr_ptr - ref_count_w;
                `uvm_info("PKT_DROP_DEBUG", $sformatf("Time=%0t: Packet drop: wr_ptr %0d -> %0d (count_w=%0d)", 
                         $time, ref_wr_ptr, ref_wr_ptr_next, ref_count_w), UVM_LOW)
            end
            
            // CRITICAL DEBUG: Track buffer writes when wr_lvl = 0
            if (ref_wr_lvl == 0) begin
                `uvm_info("BUFFER_WRITE_DEBUG", $sformatf("Time=%0t: WRITING TO BUFFER[0]: wr_en=%0b, buffer_full=%0b, state=%0d, data=0x%0h", 
                         $time, ref_wr_en, ref_buffer_full, write_state, ref_wr_data_r1), UVM_LOW)
            end
        end
        
        // Read operations using CURRENT pipeline register values (matching RTL exactly)
        // RTL uses deq_req_r (current pipeline register value) to generate rd_en, so scoreboard must do the same
        // This prevents the 1-cycle timing mismatch where rd_data_o is read even when deq_req=0
        // CRITICAL FIX: Handle concurrent read/write operations properly
        // This fixes the issue where rd_data_expected was one cycle slower than DUT in concurrent test
        // The key insight: data is available if there's data in the buffer OR if we're about to write data
        // We check for write to current read location (not concurrent read/write) to avoid negative wr_lvl
        if (ref_deq_req_r && (read_state == READ_HEADER || read_state == READ_DATA)) begin
            // Check if data is available for reading
            bit data_available = 0;
            
            if (!ref_buffer_empty) begin
                // Normal case: data available in buffer
                data_available = 1;
            end else if (ref_wr_en && (ref_wr_ptr == ref_rd_ptr)) begin
                // Special case: writing to current read location, data will be available after write
                // This ensures we don't read stale data, but also don't create negative wr_lvl
                data_available = 1;
                `uvm_info("RD_DATA_DEBUG", $sformatf("Time=%0t: WRITE to current read location: wr_ptr=%0d, rd_ptr=%0d, data will be available after write", 
                         $time, ref_wr_ptr, ref_rd_ptr), UVM_LOW)
            end
            
            if (data_available) begin
                // CRITICAL FIX: Simplified pointer-based timing - read immediately, advance pointer with delay
                // Read data directly from buffer using current pointer (immediate)
                ref_rd_data_o = ref_buffer[ref_rd_ptr[13:0]];
                // Calculate next read pointer position (will be updated on next cycle)
                ref_rd_ptr_next = ref_rd_ptr + 1;
                `uvm_info("RD_DATA_DEBUG", $sformatf("Time=%0t: Read operation: deq_req_r=%0b, state=%0d, rd_data=0x%0h, current_ptr=%0d, next_ptr=%0d (pointer advances next cycle)", 
                         $time, ref_deq_req_r, read_state, ref_rd_data_o, ref_rd_ptr, ref_rd_ptr_next), UVM_LOW)
            end else begin
                // No data available - keep pointer unchanged
                ref_rd_ptr_next = ref_rd_ptr;
                `uvm_info("RD_DATA_DEBUG", $sformatf("Time=%0t: No data available for read: deq_req_r=%0b, state=%0d, wr_en=%0b, rd_en=%0b, wr_ptr=%0d, rd_ptr=%0d, buffer_empty=%0b", 
                         $time, ref_deq_req_r, read_state, ref_wr_en, ref_rd_en, ref_wr_ptr, ref_rd_ptr, ref_buffer_empty), UVM_LOW)
            end
        end else begin
            // No read operation this cycle - keep pointer unchanged
            ref_rd_ptr_next = ref_rd_ptr;
        end
            
        // Packet length read aligns with deq_req_r in READ_HEADER (matching RTL exactly)
        if (read_state == READ_HEADER && ref_deq_req_r) begin
            ref_packet_length = ref_pck_len_buffer[ref_pck_len_rd_ptr[4:0]];
            ref_pck_len_rd_ptr = ref_pck_len_rd_ptr + 1;
            `uvm_info("PKT_LEN_READ_DEBUG", $sformatf("Time=%0t: Packet length read: deq_req_r=%0b, pck_len=%0d, ptr=%0d", 
                     $time, ref_deq_req_r, ref_packet_length, ref_pck_len_rd_ptr-1), UVM_LOW)
        end
        
        // CRITICAL FIX: Reset count_w when packet completes normally (matching RTL exactly)
        // RTL resets count_w when: (in_eop_r1 && present_state_w == WRITE_DATA) || packet_drop
        if (ref_in_eop_r1 && (write_state == WRITE_DATA)) begin
            `uvm_info("COUNT_W_DEBUG", $sformatf("Time=%0t: Packet completed normally: resetting count_w from %0d to 0 (in_eop_r1=%0b, state=%0d)", 
                     $time, ref_count_w, ref_in_eop_r1, write_state), UVM_LOW)
            ref_count_w_next = 0;
        end
        
    
        // ============================================================================
        // PHASE 9: Update previous-cycle trackers (for next cycle use)
        // ============================================================================
        ref_rd_en_prev = ref_rd_en;
        ref_wr_en_prev = ref_wr_en;
        // ref_buffer_full_prev2 = ref_buffer_full_prev;  // Two-cycle delay for overflow
        // ref_buffer_full_prev  = ref_buffer_full;
        // ref_buffer_empty_prev = ref_buffer_empty;
        // ref_overflow_prev = ref_overflow;
        ref_deq_req_prev2 = ref_deq_req_prev;
        ref_deq_req_prev = ref_deq_req_r;
        
        // Debug buffer_full timing for overflow detection
        if (ref_buffer_full != ref_buffer_full_prev) begin
            `uvm_info("BUFFER_FULL_TIMING", $sformatf("Time=%0t: buffer_full changed: %0b -> %0b (prev2=%0b for overflow)", 
                     $time, ref_buffer_full_prev, ref_buffer_full, ref_buffer_full_prev2), UVM_LOW)
        end
        
        // ============================================================================
        // PHASE 10: Update overflow/underflow detection (uses previous cycle values)
        // ============================================================================
        update_overflow_underflow(tr);             // Sets ref_pck_proc_overflow, ref_pck_proc_underflow
        
        // ============================================================================
        // PHASE 11: Update packet drop logic and outputs (moved here as requested)
        // ============================================================================
        update_packet_drop_logic(tr);              // Sets ref_packet_drop (moved to after buffer operations)
        
        // CRITICAL FIX: Recompute FSM next states after packet drop logic is calculated
        // This ensures FSM can use the correct ref_packet_drop value for state transitions
        compute_write_next_state(tr);              // Recompute write_state_next with updated ref_packet_drop
        compute_read_next_state(tr);               // Recompute read_state_next with updated ref_packet_drop
        

         // CRITICAL FIX: Calculate wr_lvl_next based on enable signals (matching RTL exactly)
        // This ensures correct wr_lvl behavior for concurrent read/write operations
        if (ref_wr_en && ref_rd_en) begin
            // Concurrent read/write: wr_lvl stays constant (both pointers advance)
            ref_wr_lvl_next = ref_wr_ptr_next - ref_rd_ptr_next - 1;
            `uvm_info("WR_LVL_NEXT", $sformatf("Time=%0t: CONCURRENT R/W: wr_lvl_next=%0d (wr_ptr_next=%0d - rd_ptr_next=%0d - 1)", 
                     $time, ref_wr_lvl_next, ref_wr_ptr_next, ref_rd_ptr_next), UVM_LOW)
        end else if (ref_wr_en) begin
            // Write only: wr_lvl increases by 1 (wr_ptr advances, rd_ptr stays)
            ref_wr_lvl_next = ref_wr_ptr_next - ref_rd_ptr_next;
            `uvm_info("WR_LVL_NEXT", $sformatf("Time=%0t: WRITE ONLY: wr_lvl_next=%0d (wr_ptr_next=%0d - rd_ptr_next=%0d)", 
                     $time, ref_wr_lvl_next, ref_wr_ptr_next, ref_rd_ptr_next), UVM_LOW)
        end else if (ref_rd_en) begin
            // Read only: wr_lvl decreases by 1 (wr_ptr stays, rd_ptr advances)
            ref_wr_lvl_next = ref_wr_ptr_next - ref_rd_ptr_next - 1;
            `uvm_info("WR_LVL_NEXT", $sformatf("Time=%0t: READ ONLY: wr_lvl_next=%0d (wr_ptr_next=%0d - rd_ptr_next=%0d)", 
                     $time, ref_wr_lvl_next, ref_wr_ptr_next, ref_rd_ptr_next), UVM_LOW)
        end else if (tr.deq_req && (read_state_next == READ_HEADER || read_state_next == READ_DATA)) begin
            // PENDING READ: deq_req is asserted and FSM will transition to read state next cycle
            // Check if data will be available for reading
            bit data_will_be_available = 0;
            if (!ref_buffer_empty) begin
                // Normal case: data available in buffer
                data_will_be_available = 1;
            end else if (ref_wr_en && (ref_wr_ptr_next == ref_rd_ptr_next)) begin
                // Special case: writing to current read location, data will be available after write
                data_will_be_available = 1;
            end
            
            if (data_will_be_available) begin
                // wr_lvl should decrease by 1 because read will happen next cycle
                ref_wr_lvl_next = ref_wr_ptr_next - ref_rd_ptr_next - 1;
                `uvm_info("WR_LVL_NEXT", $sformatf("Time=%0t: PENDING READ: wr_lvl_next=%0d (deq_req=1, next_state=%0d, wr_ptr_next=%0d - rd_ptr_next=%0d - 1, data_available=%0b)", 
                         $time, ref_wr_lvl_next, read_state_next, ref_wr_ptr_next, ref_rd_ptr_next, data_will_be_available), UVM_LOW)
            end else begin
                // No data available - wr_lvl stays constant
                ref_wr_lvl_next = ref_wr_ptr_next - ref_rd_ptr_next;
                `uvm_info("WR_LVL_NEXT", $sformatf("Time=%0t: PENDING READ (no data): wr_lvl_next=%0d (deq_req=1, next_state=%0d, wr_ptr_next=%0d - rd_ptr_next=%0d, data_available=%0b)", 
                         $time, ref_wr_lvl_next, read_state_next, ref_wr_ptr_next, ref_rd_ptr_next, data_will_be_available), UVM_LOW)
            end
        end else begin
            // No operation: wr_lvl stays constant (both pointers stay)
            ref_wr_lvl_next = ref_wr_ptr_next - ref_rd_ptr_next;
            `uvm_info("WR_LVL_NEXT", $sformatf("Time=%0t: NO OP: wr_lvl_next=%0d (wr_ptr_next=%0d - rd_ptr_next=%0d)", 
                     $time, ref_wr_lvl_next, ref_wr_ptr_next, ref_rd_ptr_next), UVM_LOW)
        end


        // Debug next states computed after packet drop logic
        `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: Next states recomputed after packet drop - WRITE: %0d -> %0d, READ: %0d -> %0d, packet_drop=%0b", 
                 $time, write_state, write_state_next, read_state, read_state_next, ref_packet_drop), UVM_LOW)
        
        // ============================================================================
        // PHASE 12: Advance states (simultaneous update matching RTL <=)
        // ============================================================================
        if (write_state != write_state_next) begin
            `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: WRITE FSM ADVANCE: %0d -> %0d", 
                     $time, write_state, write_state_next), UVM_LOW)
        end
        if (read_state != read_state_next) begin
            `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: READ FSM ADVANCE: %0d -> %0d", 
                     $time, read_state, read_state_next), UVM_LOW)
        end
        read_state_prev = read_state;  // Store previous state before advancing
        write_state = write_state_next;
        read_state  = read_state_next;
        
        // ============================================================================
        // PHASE 13: Update pipeline registers (simultaneous update matching RTL <=)
        // ============================================================================
        `uvm_info("PIPELINE_TIMING", $sformatf("Time=%0t: Updating pipeline registers for next cycle use (matching RTL <= behavior)", $time), UVM_LOW)
        update_pipeline_registers(tr);
        
        // CRITICAL FIX: Update read pointer with 1-cycle delay to match RTL timing
        // RTL registers read pointer, so it updates one cycle after deq_req_r goes high
       // ref_rd_ptr = ref_rd_ptr_next;
        // `uvm_info("RD_PTR_TIMING", $sformatf("Time=%0t: Updated rd_ptr=%0d from rd_ptr_next (1-cycle delay matching RTL)", 
        //          $time, ref_rd_ptr), UVM_LOW)
        
        // ============================================================================
        // PHASE 14: Update outputs (AFTER pipeline registers are updated)
        // ============================================================================
        update_outputs(tr);                        // Sets ref_out_sop, ref_out_eop, ref_count_r (now uses updated ref_deq_req_r)
        
        // ============================================================================
        // PHASE 15: Final updates for next cycle
        // ============================================================================
        ref_count_w_prev = ref_count_w;
        ref_count_w2_prev = ref_count_w2;  // CRITICAL FIX: Add count_w2_prev update for new RTL
        
        // CRITICAL FIX: Update count_r to match RTL's always_ff behavior
        // RTL priority: out_eop reset FIRST, then increment (matching RTL exactly)
        if (ref_out_eop) begin
            // FIRST PRIORITY: Reset count_r when out_eop is asserted (matching RTL)
            ref_count_r = 0;
            `uvm_info("COUNT_R_UPDATE", $sformatf("Time=%0t: count_r reset to 0 (out_eop=%0b) - FIRST PRIORITY", 
                     $time, ref_out_eop), UVM_LOW)
        end else if (ref_deq_req_r && (read_state_prev == READ_HEADER || read_state_prev == READ_DATA)) begin
            // SECOND PRIORITY: Increment count_r only if NOT out_eop (matching RTL)
            ref_count_r = ref_count_r + 1;
            `uvm_info("COUNT_R_UPDATE", $sformatf("Time=%0t: count_r incremented to %0d (deq_req_r=%0b, prev_state=%0d) - SECOND PRIORITY", 
                     $time, ref_count_r, ref_deq_req_r, read_state_prev), UVM_LOW)
        end
        
        // Debug count_w tracking for packet drop
        if (ref_count_w != ref_count_w_prev) begin
            `uvm_info("COUNT_W_TRACKING", $sformatf("Time=%0t: count_w changed: prev=%0d -> curr=%0d (for next cycle packet drop)", 
                     $time, ref_count_w_prev, ref_count_w), UVM_LOW)
        end
        
        // Debug count_w2 tracking for packet drop
        if (ref_count_w2 != ref_count_w2_prev) begin
            `uvm_info("COUNT_W2_TRACKING", $sformatf("Time=%0t: count_w2 changed: prev=%0d -> curr=%0d (for next cycle packet drop)", 
                     $time, ref_count_w2_prev, ref_count_w2), UVM_LOW)
        end
        
        // // ============================================================================
        // // PHASE 16: Buffer synchronization
        // // ============================================================================
        // // CRITICAL FIX: Update pointers for next cycle (matching RTL always_ff behavior)
        // ref_wr_ptr = ref_wr_ptr_next;  // Update write pointer
        // ref_rd_ptr = ref_rd_ptr_next;  // Update read pointer
        
        // // CRITICAL FIX: Calculate wr_lvl based on pointers (matching RTL exactly)
        // // RTL: wr_lvl = wr_ptr - rd_ptr
        // ref_wr_lvl = ref_wr_ptr - ref_rd_ptr;

        // update_buffer_states();
        
        // CRITICAL FIX: Reset read pointer when wr_lvl is reset to 0 (buffer empty)
        // This ensures read pointer stays synchronized with write level
        if (ref_wr_lvl == 0 && ref_rd_ptr != 0) begin
            `uvm_info("BUFFER_SYNC_DEBUG", $sformatf("Time=%0t: Buffer empty: resetting read pointer from %0d to 0 (wr_lvl=%0d)", 
                     $time, ref_rd_ptr, ref_wr_lvl), UVM_LOW)
            ref_rd_ptr = 0;
        end
        
        // ============================================================================
        // PHASE 17: DEBUG - Final state verification
        // ============================================================================
        // Debug state alignment for write enable generation
        `uvm_info("STATE_ALIGNMENT", $sformatf("Time=%0t: State alignment - Scoreboard write_state=%0d, DUT present_state=%0d, ref_wr_en=%0b, enq_req_r=%0b, enq_req_curr=%0b", 
                 $time, write_state, tr.pck_proc_int_mem_fsm_rstn ? 0 : 2, ref_wr_en, ref_enq_req_r, tr.enq_req), UVM_LOW)
        
        // Additional debug: Show when registered enq_req is used
        if (ref_enq_req_r != tr.enq_req) begin
            `uvm_info("ENQ_REQ_TIMING", $sformatf("Time=%0t: enq_req changed: registered=%0b -> curr=%0b, using registered for wr_en=%0b", 
                     $time, ref_enq_req_r, tr.enq_req, ref_wr_en), UVM_LOW)
        end
        
        // Additional debug: Show the exact timing relationship
        `uvm_info("TIMING_DEBUG", $sformatf("Time=%0t: Timing - enq_req_curr=%0b, enq_req_r=%0b, enq_req_r1=%0b, wr_en=%0b, write_state=%0d", 
                 $time, tr.enq_req, ref_enq_req_r, ref_enq_req_r1, ref_wr_en, write_state), UVM_LOW)
        
        // Enhanced debug wr_lvl calculation with more details
        `uvm_info("WR_LVL_DEBUG", $sformatf("Time=%0t: wr_lvl_next calc: wr_en=%0b, rd_en=%0b, buffer_full=%0b, buffer_empty=%0b, wr_lvl_next=%0d, current_wr_lvl=%0d, packet_drop=%0b, count_w=%0d", 
                 $time, ref_wr_en, ref_rd_en, ref_buffer_full, ref_buffer_empty, ref_wr_lvl_next, ref_wr_lvl, ref_packet_drop, ref_count_w), UVM_LOW)
        
        // Additional debug: Track when write level should change
        if (ref_wr_lvl_next != ref_wr_lvl) begin
            `uvm_info("WR_LVL_CHANGE", $sformatf("Time=%0t: WR_LVL CHANGE DETECTED: %0d -> %0d (wr_en=%0b, rd_en=%0b, packet_drop=%0b)", 
                     $time, ref_wr_lvl, ref_wr_lvl_next, ref_wr_en, ref_rd_en, ref_packet_drop), UVM_LOW)
        end
        
        // CRITICAL FIX: ref_wr_lvl is NOT updated here - it's updated in write() after comparison
        // This ensures comparison uses current cycle value, but wr_lvl is ready for next cycle
        // This matches RTL where wr_lvl updates at clock edge for next cycle use
    endfunction

    function void handle_reset_logic(pkt_proc_seq_item tr);
        // Asynchronous active-low reset (highest priority)
        if (!tr.pck_proc_int_mem_fsm_rstn) begin
            `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: ASYNC RESET: Resetting all states to IDLE", $time), UVM_LOW)
            // Set reset active flag (matching DUT async reset behavior)
            ref_reset_active = 1;
            
            // Reset all state machines and registers
            write_state = IDLE_W;
            read_state = IDLE_R;
            
            // Reset pointers and counters
            ref_wr_ptr = 0;           // Reset write pointer
            ref_wr_ptr_next = 0;      // Reset next write pointer
            ref_rd_ptr = 0;
            ref_rd_ptr_next = 0;  // Reset next cycle's read pointer
            ref_pck_len_wr_ptr = 0;
            ref_pck_len_rd_ptr = 0;
            ref_wr_lvl = 0;
            ref_count_w_next = 0;       // Set next count_w to 0
            ref_count_w = 0;
            ref_count_w_prev = 0;       // Initialize previous count_w
            ref_count_w2 = 0;           // Second count_w starts at 0
            ref_count_w2_next = 0;      // Next count_w2 starts at 0
            ref_count_w2_prev = 0;      // Initialize previous count_w2
            ref_count_r = 0;
            ref_packet_length = 0;
            ref_packet_length_w = 0;
            `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: ref_packet_length_w reset to 0 (ASYNC RESET)", $time), UVM_LOW)
            
            // Reset buffer states
            //ref_buffer_full = 0;
            //ref_buffer_empty = 1;
            ref_pck_len_full = 0;
            ref_pck_len_empty = 1;
            
            // Reset flags
            ref_pck_proc_overflow = 0;
            ref_pck_proc_underflow = 0;
            ref_packet_drop = 0;
            ref_packet_drop_prev = 0;
            invalid_1 = 0;
            invalid_3 = 0;
            invalid_4 = 0;
            invalid_5 = 0;
            invalid_6 = 0;
            any_invalid_condition = 0;
            ref_overflow = 0;
            
            // Reset outputs
            ref_out_sop = 0;
            ref_out_eop = 0;
            ref_rd_data_o = 0;
            //ref_pck_proc_almost_full = 0;
            //ref_pck_proc_almost_empty = 0;
            
            // Reset pipeline registers
            ref_in_sop_r = 0; ref_in_sop_r1 = 0; ref_in_sop_r2 = 0;
            ref_in_eop_r = 0; ref_in_eop_r1 = 0; ref_in_eop_r2 = 0;
            ref_enq_req_r = 0; ref_enq_req_r1 = 0;
            ref_wr_data_r = 0; ref_wr_data_r1 = 0;
            ref_pck_len_valid_r = 0; ref_pck_len_valid_r1 = 0;
            ref_pck_len_i_r = 0; ref_pck_len_i_r1 = 0;
            ref_deq_req_r = 0;
            
            // Reset additional signals
            ref_empty_de_assert = 0;
            ref_buffer_empty_r = 1;
            ref_wr_en = 0;
            ref_rd_en = 0;
            ref_wr_lvl_next = 0;
            
            return; // Exit early - no further processing during reset
        end
        
        // Check if reset was just de-asserted (transition from reset to normal operation)
        if (ref_reset_active && tr.pck_proc_int_mem_fsm_rstn) begin
            `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: RESET DE-ASSERTED: Returning to normal operation", $time), UVM_LOW)
            ref_reset_active = 0;
        end
        
        // Synchronous active-high software reset (second priority)
        if (tr.pck_proc_int_mem_fsm_sw_rstn) begin
            `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: SYNC RESET: Resetting all states to IDLE", $time), UVM_LOW)
            // Set reset active flag for software reset
            ref_reset_active = 1;
            
            // Reset all state machines and registers
            write_state = IDLE_W;
            read_state = IDLE_R;
            
            // Reset pointers and counters
            ref_wr_ptr = 0;           // Reset write pointer
            ref_wr_ptr_next = 0;      // Reset next write pointer
            ref_rd_ptr = 0;
            ref_rd_ptr_next = 0;  // Reset next cycle's read pointer
            ref_pck_len_wr_ptr = 0;
            ref_pck_len_rd_ptr = 0;
            ref_wr_lvl = 0;
            ref_count_w = 0;       // Set next count_w to 0
            ref_count_w_next = 0;       // Set next count_w to 0
            ref_count_w_prev = 0;       // Initialize previous count_w
            ref_count_w2 = 0;           // Second count_w starts at 0
            ref_count_w2_next = 0;      // Next count_w2 starts at 0
            ref_count_w2_prev = 0;      // Initialize previous count_w2
            ref_count_r = 0;
            ref_packet_length = 0;
            ref_packet_length_w = 0;
            `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: ref_packet_length_w reset to 0 (SYNC RESET)", $time), UVM_LOW)
            
            // Reset buffer states
            //ref_buffer_full = 0;
            //ref_buffer_empty = 1;
            ref_pck_len_full = 0;
            ref_pck_len_empty = 1;
            
            // Reset flags
            ref_pck_proc_overflow = 0;
            ref_pck_proc_underflow = 0;
            ref_packet_drop = 0;
            ref_packet_drop_prev = 0;
            invalid_1 = 0;
            invalid_3 = 0;
            invalid_4 = 0;
            invalid_5 = 0;
            invalid_6 = 0;
            any_invalid_condition = 0;
            ref_overflow = 0;
            
            // Reset outputs
            ref_out_sop = 0;
            ref_out_eop = 0;
            ref_rd_data_o = 0;
            //ref_pck_proc_almost_full = 0;
            //ref_pck_proc_almost_empty = 0;
            
            // Reset pipeline registers
            ref_in_sop_r = 0; ref_in_sop_r1 = 0; ref_in_sop_r2 = 0;
            ref_in_eop_r = 0; ref_in_eop_r1 = 0; ref_in_eop_r2 = 0;
            ref_enq_req_r = 0; ref_enq_req_r1 = 0;
            ref_wr_data_r = 0; ref_wr_data_r1 = 0;
            ref_pck_len_valid_r = 0; ref_pck_len_valid_r1 = 0;
            ref_pck_len_i_r = 0; ref_pck_len_i_r1 = 0;
            ref_deq_req_r = 0;
            
            // Reset additional signals
            ref_empty_de_assert = 0;
            ref_buffer_empty_r = 1;
            ref_wr_en = 0;
            ref_rd_en = 0;
            ref_wr_lvl_next = 0;
            ref_rd_ptr_next = 0;  // Reset next cycle's read pointer

            data_available = 0;
            data_available_next = 0;
            data_available_for_comparison = 0;
            
            return; // Exit early - no further processing during reset
        end
        
        // Check if software reset was just de-asserted
        if (ref_reset_active && !tr.pck_proc_int_mem_fsm_sw_rstn) begin
            `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: SOFTWARE RESET DE-ASSERTED: Returning to normal operation", $time), UVM_LOW)
            ref_reset_active = 0;
        end
    endfunction

    function void update_pipeline_registers(pkt_proc_seq_item tr);
        // Pipeline registers (matching RTL exactly)
        // CRITICAL FIX: Correct pipeline order - shift values from previous cycle
        ref_in_sop_r2 = ref_in_sop_r1;  // 2-cycle delayed in_sop
        ref_in_sop_r1 = ref_in_sop_r;   // 1-cycle delayed in_sop  
        ref_in_sop_r = tr.in_sop;       // Current cycle in_sop
        
        ref_in_eop_r2 = ref_in_eop_r1;  // 2-cycle delayed in_eop
        ref_in_eop_r1 = ref_in_eop_r;   // 1-cycle delayed in_eop
        ref_in_eop_r = tr.in_eop;       // Current cycle in_eop
        
        ref_enq_req_r1 = ref_enq_req_r; // 1-cycle delayed enq_req
        ref_enq_req_r = tr.enq_req;     // Current cycle enq_req
        
        ref_wr_data_r1 = ref_wr_data_r; // 1-cycle delayed wr_data
        ref_wr_data_r = tr.wr_data_i;   // Current cycle wr_data
        
        ref_pck_len_valid_r1 = ref_pck_len_valid_r;  // 1-cycle delayed pck_len_valid
        ref_pck_len_valid_r = tr.pck_len_valid;      // Current cycle pck_len_valid
        
        ref_pck_len_i_r1 = ref_pck_len_i_r;         // 1-cycle delayed pck_len_i
        ref_pck_len_i_r = tr.pck_len_i;             // Current cycle pck_len_i
        
        // Debug pipeline register updates
        `uvm_info("PIPELINE_UPDATE", $sformatf("Time=%0t: Pipeline updated - in_sop: %0b->%0b->%0b, in_eop: %0b->%0b->%0b", 
                 $time, tr.in_sop, ref_in_sop_r1, ref_in_sop_r2, tr.in_eop, ref_in_eop_r1, ref_in_eop_r2), UVM_LOW)
        
        // Model RTL register on deq_req: stage and then register
        ref_deq_req_r1 = tr.deq_req;  // sample input
        ref_deq_req_r  = ref_deq_req_r1; // registered output (1-cycle delayed)
        ref_empty_de_assert = tr.empty_de_assert;
        
        // CRITICAL FIX: Do NOT update ref_wr_lvl here - it should update on NEXT cycle like RTL
        // The RTL wr_lvl updates on the NEXT clock edge, not the current one
        // ref_wr_lvl = ref_wr_lvl_next;  // REMOVED - this was causing 1-cycle ahead behavior
        
        // Debug write level timing
        `uvm_info("WR_LVL_TIMING", $sformatf("Time=%0t: ref_wr_lvl_next=%0d calculated, but ref_wr_lvl=%0d NOT updated yet (matching RTL always_ff timing)", 
                 $time, ref_wr_lvl_next, ref_wr_lvl), UVM_LOW)
    endfunction

    function void compute_write_next_state(pkt_proc_seq_item tr);
        unique case (write_state)
            IDLE_W: begin
                // Use current cycle values (matching RTL behavior exactly)
                if (tr.enq_req && tr.in_sop) begin
                    write_state_next = WRITE_HEADER;
                    `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: WRITE FSM: IDLE_W -> WRITE_HEADER (enq_req=%0b, in_sop=%0b)", 
                             $time, tr.enq_req, tr.in_sop), UVM_LOW)
                end else begin
                    write_state_next = IDLE_W;
                end
            end
            
            WRITE_HEADER: begin
                // Use current cycle values (matching RTL behavior exactly)
                if (tr.in_sop) begin
                    write_state_next = WRITE_HEADER;
                    `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: WRITE FSM: WRITE_HEADER -> WRITE_HEADER (in_sop=%0b)", 
                             $time, tr.in_sop), UVM_LOW)
                end else if (ref_packet_drop) begin
                    // CRITICAL FIX: When packet drop is detected, go to IDLE_W instead of ERROR
                    // This matches RTL behavior where invalid packets are dropped and FSM returns to idle
                    write_state_next = IDLE_W;
                    `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: WRITE FSM: WRITE_HEADER -> IDLE_W (packet_drop=%0b, invalid packet dropped)", 
                             $time, ref_packet_drop), UVM_LOW)
                    
                    // CRITICAL DEBUG: Show why packet drop occurred
                    if (invalid_1) begin
                        `uvm_info("STATE_TRANSITION_DEBUG", $sformatf("Time=%0t: Transitioning to IDLE_W due to invalid_1: in_sop_r1=%0b && in_eop_r1=%0b (same cycle)", 
                                 $time, ref_in_sop_r1, ref_in_eop_r1), UVM_LOW)
                    end
                end else begin
                    write_state_next = WRITE_DATA;
                    `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: WRITE FSM: WRITE_HEADER -> WRITE_DATA (advance to data)", $time), UVM_LOW)
                end
            end
            
            WRITE_DATA: begin
                // CRITICAL FIX: Check for packet drop in WRITE_DATA state as well
                if (ref_packet_drop) begin
                    // When packet drop is detected in WRITE_DATA, go to IDLE_W
                    write_state_next = IDLE_W;
                    `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: WRITE FSM: WRITE_DATA -> IDLE_W (packet_drop=%0b, invalid packet dropped)", 
                             $time, ref_packet_drop), UVM_LOW)
                    
                    // CRITICAL DEBUG: Show why packet drop occurred
                    if (invalid_3 || invalid_4 || invalid_5 || invalid_6) begin
                        `uvm_info("STATE_TRANSITION_DEBUG", $sformatf("Time=%0t: Transitioning to IDLE_W due to invalid_3 || invalid_4 || invalid_5 || invalid_6", 
                                 $time), UVM_LOW)
                    end
                end else if ((tr.in_sop && ref_in_eop_r1 && tr.enq_req) || (tr.in_sop && tr.enq_req)) begin
                    write_state_next = WRITE_HEADER;
                    `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: WRITE FSM: WRITE_DATA -> WRITE_HEADER (next_data_ready: in_sop=%0b, in_eop_r1=%0b, enq_req=%0b)", 
                             $time, tr.in_sop, ref_in_eop_r1, tr.enq_req), UVM_LOW)
                end else if (ref_in_eop_r1 && !tr.in_sop && !tr.enq_req) begin
                    write_state_next = IDLE_W;
                    `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: WRITE FSM: WRITE_DATA -> IDLE_W (next_data_nt_ready: in_eop_r1=%0b, in_sop=%0b, enq_req=%0b)", 
                             $time, ref_in_eop_r1, tr.in_sop, tr.enq_req), UVM_LOW)
                end else begin
                    write_state_next = WRITE_DATA;
                end
            end
            
            default: begin
                write_state_next = IDLE_W;
                `uvm_error("STATE_TRANSITION", $sformatf("Time=%0t: WRITE FSM: Unknown state %0d, resetting to IDLE_W", $time, write_state))
            end
        endcase
    endfunction

    function void compute_read_next_state(pkt_proc_seq_item tr);
        // CRITICAL FIX: Read state machine now properly handles write to current read location
        // When wr_ptr == rd_ptr and wr_en is high, data will be available after write
        // This prevents the 1-cycle delay in read operations that was causing rd_data_expected mismatch
        unique case (read_state)
            IDLE_R: begin
                // Use registered values (matching RTL behavior exactly)
                // CRITICAL FIX: Handle concurrent read/write operations properly
                data_available = 0;
                if (!ref_buffer_empty) begin
                    // Normal case: data available in buffer
                    data_available = 1;
                end else if (ref_wr_en && (ref_wr_ptr == ref_rd_ptr)) begin
                    // Special case: writing to current read location, data will be available after write
                    data_available = 1;
                end
                
                if (ref_deq_req_r && data_available) begin
                    read_state_next = READ_HEADER;
                    `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: READ FSM: IDLE_R -> READ_HEADER (deq_req_r=%0b, data_available=%0b, wr_en=%0b, rd_en=%0b, wr_ptr=%0d, rd_ptr=%0d)", 
                             $time, ref_deq_req_r, data_available, ref_wr_en, ref_rd_en, ref_wr_ptr, ref_rd_ptr), UVM_LOW)
                end else begin
                    read_state_next = IDLE_R;
                end
            end
            
            READ_HEADER: begin
                read_state_next = READ_DATA;
                `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: READ FSM: READ_HEADER -> READ_DATA (advance to data)", $time), UVM_LOW)
            end
            
            READ_DATA: begin
                // CRITICAL FIX: Handle concurrent read/write operations properly
                data_available = 0;
                if (!ref_buffer_empty) begin
                    // Normal case: data available in buffer
                    data_available = 1;
                end else if (ref_wr_en && (ref_wr_ptr == ref_rd_ptr)) begin
                    // Special case: writing to current read location, data will be available after write
                    data_available = 1;
                end
                
                if (!data_available) begin
                    read_state_next = IDLE_R;
                    `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: READ FSM: READ_DATA -> IDLE_R (no data available - wr_en=%0b, rd_en=%0b, wr_ptr=%0d, rd_ptr=%0d, buffer_empty=%0b)", 
                             $time, ref_wr_en, ref_rd_en, ref_wr_ptr, ref_rd_ptr, ref_buffer_empty), UVM_LOW)
                end else if ((ref_count_r == (ref_packet_length - 1)) && ref_deq_req_r && data_available) begin
                    read_state_next = READ_HEADER;  // Next packet
                    `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: READ FSM: READ_DATA -> READ_HEADER (next packet: count_r=%0d, pck_len=%0d, deq_req_r=%0b)", 
                             $time, ref_count_r, ref_packet_length, ref_deq_req_r), UVM_LOW)
                end else if ((ref_count_r == (ref_packet_length - 1)) && (!ref_deq_req_r || !data_available)) begin
                    read_state_next = IDLE_R;  // End of packet
                    `uvm_info("STATE_TRANSITION", $sformatf("Time=%0t: READ FSM: READ_DATA -> IDLE_R (end of packet: count_r=%0d, pck_len=%0d, deq_req_r=%0b)", 
                             $time, ref_count_r, ref_packet_length, ref_deq_req_r), UVM_LOW)
                end else begin
                    read_state_next = READ_DATA;  // Continue reading
                end
            end
        endcase
    endfunction

    function void generate_write_read_enables(pkt_proc_seq_item tr);
        // CRITICAL FIX: Update to match new RTL behavior
        // New RTL sets wr_en=1 when pck_invalid=1 (packet_drop=1) to write the invalid packet data
        if (ref_packet_drop) begin
            ref_wr_en = 1;  // Write invalid packet data (matching new RTL behavior)
            `uvm_info("WR_EN_DEBUG", $sformatf("Time=%0t: Packet drop detected - setting wr_en=1 to write invalid packet data (new RTL behavior)", $time), UVM_LOW)
            
            // CRITICAL DEBUG: Show buffer state when packet drop triggers write
            `uvm_info("WR_EN_DEBUG", $sformatf("Time=%0t: Buffer state during packet drop: wr_lvl=%0d, count_w=%0d, state=%0d", 
                     $time, ref_wr_lvl, ref_count_w, write_state), UVM_LOW)
        end else begin
            // CRITICAL FIX: Use ref_enq_req_r (1-cycle delayed) to match RTL exactly
            // RTL uses enq_req_r (1-cycle delayed enq_req) for wr_en generation
            case (write_state)
                IDLE_W: begin
                    ref_wr_en = 0;
                end
                WRITE_HEADER: begin
                    // RTL: wr_en = (enq_req_r) ? 1 : 0
                    ref_wr_en = (ref_enq_req_r) ? 1 : 0;
                end
                WRITE_DATA: begin
                    // RTL: wr_en = (enq_req_r) ? 1 : 0
                    ref_wr_en = (ref_enq_req_r) ? 1 : 0;
                end
                default: begin
                    ref_wr_en = 0;
                end
            endcase
        end
        
        // Read enable logic (unchanged)
        case (read_state)
            IDLE_R: begin
                ref_rd_en = 0;
            end
            READ_HEADER: begin
                ref_rd_en = (tr.deq_req) ? 1 : 0;
            end
            READ_DATA: begin
                ref_rd_en = (tr.deq_req) ? 1 : 0;
            end
            default: begin
                ref_rd_en = 0;
            end
        endcase
        
        `uvm_info("WR_RD_EN_DEBUG", $sformatf("Time=%0t: Generated - wr_en=%0b (packet_drop=%0b, state=%0d, enq_req_r=%0b, enq_req_curr=%0b), rd_en=%0b (state=%0d, deq_req=%0b)", 
                 $time, ref_wr_en, ref_packet_drop, write_state, ref_enq_req_r, tr.enq_req, ref_rd_en, read_state, tr.deq_req), UVM_LOW)
    endfunction

    function void update_packet_drop_logic(pkt_proc_seq_item tr);
         // CRITICAL: Reset packet_drop to 0 EVERY cycle (matching RTL always_comb)
          ref_packet_drop = 0;  // Default value every cycle
        
        // Calculate packet drop logic (matching RTL exactly)
        // pck_invalid = (invalid_1 || invalid_3 || invalid_4 || invalid_5 || invalid_6) && enq_req
        // invalid_1 = in_sop && in_eop
        // invalid_3 = in_sop && (~in_eop_r1) && (write_state == WRITE_DATA)
        // invalid_4 = (count_w < (packet_length_w - 1)) && (packet_length_w != 0) && (in_eop_r1)
        // invalid_5 = ((count_w == (packet_length_w - 1)) || (packet_length_w == 0)) && (~in_eop_r1) && (write_state == WRITE_DATA)
        // invalid_6 = pck_proc_overflow

        // Use WRITE-PATH packet length for these checks
        // CRITICAL FIX: Use registered values for invalid_1 to match DUT timing
        // DUT has registered versions of in_sop and in_eop, so invalid_1 should use _r1 values
        invalid_1 = (ref_in_sop_r1 && ref_in_eop_r1);
        
        // CRITICAL DEBUG: Show when invalid_1 is detected (in_sop and in_eop at same time)
        if (invalid_1) begin
            `uvm_info("INVALID_1_DETECTION", $sformatf("Time=%0t: INVALID_1 DETECTED: in_sop_r1=%0b && in_eop_r1=%0b (same cycle), current_state=%0d, should transition to IDLE_W", 
                     $time, ref_in_sop_r1, ref_in_eop_r1, write_state), UVM_LOW)
        end
        
        invalid_3 = (ref_in_sop_r1 && (~ref_in_eop_r1) && (write_state == WRITE_HEADER));
        // CRITICAL FIX: RTL uses current count_w but registered in_eop_r1 for invalid_4
        // invalid_4 = (count_w < (pck_len_r2 - 1)) && (pck_len_r2 != 0) && (in_eop_r1)
        invalid_4 = (write_state == WRITE_DATA) && 
                        ((ref_count_w < (ref_packet_length_w - 1)) && (ref_packet_length_w != 0) && (ref_in_eop_r1));
        // CRITICAL FIX: RTL uses current count_w but registered in_eop_r1 for invalid_5
        // invalid_5 = ((count_w == pck_len_r2-1) || (pck_len_r2 == 0)) && (~in_eop_r1) && (present_state_w==WRITE_DATA)
        // RTL uses pck_len_r2 (registered packet length) and in_eop_r1 (registered in_eop)
        invalid_5 = (((ref_count_w == (ref_packet_length_w - 1)) && (ref_packet_length_w != 0)) && (~ref_in_eop_r1) && (write_state == WRITE_DATA));
        // CRITICAL FIX: invalid_6 should detect overflow immediately when buffer is full and write is attempted
        // This ensures pck_invalid is detected in the same cycle as the DUT, without circular dependency
        // invalid_6 = (enq_req && buffer_full) - immediate overflow detection
        // NOTE: Use current cycle buffer_full for immediate detection, not delayed version
        invalid_6 = (tr.enq_req && ref_buffer_full);

        // CRITICAL FIX: Track invalid conditions across cycles to match DUT behavior
        // The DUT's pck_invalid requires both invalid condition AND enq_req, but the timing might be different
        // We need to detect invalid conditions and then assert packet_drop when enq_req is high
        any_invalid_condition = (invalid_1 || invalid_3 || invalid_4 || invalid_5 || invalid_6);
        
        // Debug: Show condition calculations that use ref_packet_length_w
        `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: invalid_1=%0b (in_sop_r1=%0b && in_eop_r1=%0b), invalid_3=%0b (ref_in_sop_r1=%0b && ~ref_in_eop_r1=%0b && state=%0d)", 
                 $time, invalid_1, ref_in_sop_r1, ref_in_eop_r1, invalid_3, ref_in_sop_r1, ref_in_eop_r1, write_state), UVM_LOW)
        `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: invalid_4=%0b (count_w=%0d < pck_len_w-1=%0d && pck_len_w!=0=%0b && ref_in_eop_r1=%0b), invalid_5=%0b (count_w=%0d == pck_len_w-1=%0d || pck_len_w==0=%0b && ~in_eop_r1=%0b && state=%0d), invalid_6=%0b (overflow=%0b)", 
                 $time, invalid_4, ref_count_w, ref_packet_length_w-1, (ref_packet_length_w != 0), ref_in_eop_r1, invalid_5, ref_count_w, ref_packet_length_w-1, (ref_packet_length_w == 0), ref_in_eop_r1, write_state, invalid_6, ref_pck_proc_overflow), UVM_LOW)

        // CRITICAL FIX: RTL emulation - Use DUT's packet_drop signal directly (matching RTL exactly)
        // RTL generates packet_drop as a combinational output based on pck_invalid logic
        // Scoreboard should use the DUT's packet_drop signal to match RTL behavior exactly
        if (tr.packet_drop) begin
            // DUT detected packet drop - verify our logic matches
            if (any_invalid_condition && tr.enq_req) begin
                `uvm_info("PKT_DROP_DEBUG", $sformatf("Time=%0t: DUT packet_drop=1 confirmed: enq_req=1, state=%0d, invalid_1=%0b, invalid_3=%0b, invalid_4=%0b", 
                         $time, write_state, invalid_1, invalid_3, invalid_4), UVM_LOW)
                `uvm_info("PKT_DROP_DEBUG", $sformatf("Time=%0t: invalid_5=%0b, invalid_6=%0b, count_w=%0d, pck_len_w=%0d, in_sop_r1=%0b, in_eop_r1=%0b", 
                         $time, invalid_5, invalid_6, ref_count_w, ref_packet_length_w, ref_in_sop_r1, ref_in_eop_r1), UVM_LOW)
                
                // Additional debug for invalid_1 specifically
                if (invalid_1) begin
                    `uvm_info("INVALID_1_DEBUG", $sformatf("Time=%0t: INVALID_1 triggered: in_sop_r1=%0b && in_eop_r1=%0b", 
                             $time, ref_in_sop_r1, ref_in_eop_r1), UVM_LOW)
                end

                // Additional debug for invalid_3 specifically
                if (invalid_3) begin
                    `uvm_info("INVALID_3_DEBUG", $sformatf("Time=%0t: INVALID_3 triggered: in_sop=%0b && ~in_eop_r1=%0b && state=%0d", 
                             $time, tr.in_sop, ref_in_eop_r1, write_state), UVM_LOW)
                end
                
                // Additional debug for invalid_4 specifically
                if (invalid_4) begin
                    `uvm_info("INVALID_4_DEBUG", $sformatf("Time=%0t: INVALID_4 triggered: state=%0d, count_w=%0d < (pck_len_w-1)=%0d && pck_len_w!=0=%0b && in_eop_r1=%0b", 
                             $time, write_state, ref_count_w, ref_packet_length_w-1, (ref_packet_length_w != 0), ref_in_eop_r1), UVM_LOW)
                end
                
                // Additional debug for invalid_5 specifically
                if (invalid_5) begin
                    `uvm_info("INVALID_5_DEBUG", $sformatf("Time=%0t: INVALID_5 triggered: count_w=%0d == (pck_len_w-1)=%0d || pck_len_w==0=%0b && ~in_eop_r1=%0b && state=%0d", 
                             $time, ref_count_w, ref_packet_length_w-1, (ref_packet_length_w == 0), ref_in_eop_r1, write_state), UVM_LOW)
                end
                
                // Additional debug for invalid_6 specifically
                if (invalid_6) begin
                    `uvm_info("INVALID_6_DEBUG", $sformatf("Time=%0t: INVALID_6 triggered: enq_req=%0b && buffer_full=%0b (immediate overflow detection)", 
                             $time, tr.enq_req, ref_buffer_full), UVM_LOW)
                end
                
                ref_packet_drop = 1;  // Confirm packet drop
            end else if (any_invalid_condition && !tr.enq_req) begin
                // CRITICAL FIX: If invalid condition exists but enq_req=0, still set packet_drop=1
                // This matches RTL behavior where packet_drop persists once invalid condition is detected
                `uvm_info("PKT_DROP_DEBUG", $sformatf("Time=%0t: Invalid condition detected but enq_req=0: invalid_1=%0b, invalid_3=%0b, invalid_4=%0b, invalid_5=%0b, invalid_6=%0b", 
                         $time, invalid_1, invalid_3, invalid_4, invalid_5, invalid_6), UVM_LOW)
                ref_packet_drop = 1;
            end else begin
                // DUT says packet_drop=1 but our logic doesn't match - this indicates a mismatch
                `uvm_warning("PKT_DROP_MISMATCH", $sformatf("Time=%0t: DUT packet_drop=1 but scoreboard logic doesn't match: enq_req=%0b, invalid_conditions=%0b, state=%0d", 
                         $time, tr.enq_req, any_invalid_condition, write_state))
                ref_packet_drop = 1;  // Use DUT's value to maintain consistency
            end
        end else begin
            // DUT says packet_drop=0 - verify our logic matches
            if (any_invalid_condition && tr.enq_req) begin
                // This indicates a potential mismatch - DUT should have detected packet drop
                `uvm_warning("PKT_DROP_MISMATCH", $sformatf("Time=%0t: Scoreboard detected invalid condition but DUT packet_drop=0: enq_req=%0b, invalid_conditions=%0b, state=%0d", 
                         $time, tr.enq_req, any_invalid_condition, write_state))
            end
            ref_packet_drop = 0;  // Use DUT's value
        end
        
        // Store previous value for next cycle
        ref_packet_drop_prev = ref_packet_drop;
    endfunction

    function void update_buffer_operations(pkt_proc_seq_item tr);
        // CRITICAL FIX: Buffer write operations moved to main function after generate_write_read_enables()
        // This ensures the first write at wr_lvl=0 uses the correct wr_en value
        
        // CRITICAL FIX: Check packet drop BEFORE performing any buffer operations
        // If packet drop is detected, skip all write operations to prevent incorrect count_w/wr_ptr increments
        if (!ref_packet_drop) begin
            // Packet length buffer operations (matching RTL exactly)
            // RTL writes to pck_len_buffer in WRITE_HEADER state regardless of wr_en
            if (write_state == WRITE_HEADER) begin
                // Use RTL logic exactly: pck_len_r2 = (pck_len_valid_r1) ? pck_len_i_r1 : ((in_sop_r1) ? wr_data_r1[11:0] : packet_length)
                // CRITICAL: These _r1 values contain the PREVIOUS cycle's values (when in_sop=1, pck_len_valid=1)
                bit [11:0] pck_len_r2_value;
                if (ref_pck_len_valid_r1) begin
                    pck_len_r2_value = ref_pck_len_i_r1;
                    `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: WRITE_HEADER: Using pck_len_i_r1=%0d (pck_len_valid_r1=1)", 
                             $time, ref_pck_len_i_r1), UVM_LOW)
                end else if (ref_in_sop_r1) begin
                    pck_len_r2_value = ref_wr_data_r1[11:0];
                    `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: WRITE_HEADER: Using wr_data_r1[11:0]=%0d (in_sop_r1=1)", 
                             $time, ref_wr_data_r1[11:0]), UVM_LOW)
                end else begin
                    pck_len_r2_value = ref_packet_length_w;  // Keep previous value
                    `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: WRITE_HEADER: Using prev_packet_length=%0d (both conditions false)", 
                             $time, ref_packet_length_w), UVM_LOW)
                end
                
                // Write to packet length buffer (matching RTL pck_len_wr_en = 1'b1 in WRITE_HEADER)
                ref_pck_len_buffer[ref_pck_len_wr_ptr[4:0]] = pck_len_r2_value;
                ref_pck_len_wr_ptr = ref_pck_len_wr_ptr + 1;
                
                // Update write-path packet length mirror for pck_invalid checks
                ref_packet_length_w = pck_len_r2_value;
                
                // Debug print for packet length assignment
                `uvm_info("PACKET_LENGTH_DEBUG", $sformatf("Time=%0t: WRITE_HEADER: pck_len_r2=%0d (pck_len_valid_r1=%0b, in_sop_r1=%0b, pck_len_i_r1=%0d, wr_data_r1[11:0]=%0d, prev_packet_length=%0d)", 
                         $time, pck_len_r2_value, ref_pck_len_valid_r1, ref_in_sop_r1, ref_pck_len_i_r1, ref_wr_data_r1[11:0], ref_packet_length_w), UVM_LOW)
            end
        end else begin
            // CRITICAL FIX: When packet drop is detected, skip all write operations
            // This prevents incorrect count_w and wr_ptr increments that would affect wr_lvl
            `uvm_info("PKT_DROP_DEBUG", $sformatf("Time=%0t: Packet drop detected - skipping buffer write operations to prevent incorrect count_w/wr_ptr increments", $time), UVM_LOW)
        end
        

        
        // CRITICAL FIX: Reset count_w when packet completes normally (matching RTL exactly)
        // RTL resets count_w when: (in_eop_r1 && present_state_w == WRITE_DATA) || packet_drop
        if (ref_in_eop_r1 && (write_state == WRITE_DATA)) begin
            `uvm_info("COUNT_W_DEBUG", $sformatf("Time=%0t: Packet completed normally: resetting count_w from %0d to 0 (in_eop_r1=%0b, state=%0d)", 
                     $time, ref_count_w, ref_in_eop_r1, write_state), UVM_LOW)
            ref_count_w_next = 0;
        end
    endfunction

    function void update_buffer_states();
        // CRITICAL FIX: Buffer full should be based on wr_lvl, not pointer comparison
        // DUT logic: pck_proc_full = 1 when wr_lvl == DEPTH (buffer is full)
        // This matches the actual RTL behavior
        ref_buffer_full = (ref_wr_lvl == DEPTH) ? 1 : 0;  // Use parameter instead of hardcoded value
        
        // CRITICAL FIX: Buffer empty should be based on wr_lvl, not pointer comparison
        // DUT logic: pck_proc_empty = 1 when wr_lvl > 0 (buffer has data)
        // This matches the actual RTL behavior
        ref_buffer_empty = (ref_wr_lvl > 0) ? 0 : 1;
        
        // CRITICAL DEBUG: Track buffer state changes, especially when wr_lvl = 0
        if (ref_wr_lvl == 0) begin
            `uvm_info("BUFFER_STATE_DEBUG", $sformatf("Time=%0t: BUFFER STATE at wr_lvl=0: full=%0b, empty=%0b, wr_en=%0b, rd_en=%0b", 
                     $time, ref_buffer_full, ref_buffer_empty, ref_wr_en, ref_rd_en), UVM_LOW)
        end
        
        // Debug buffer state
        `uvm_info("BUFFER_DEBUG", $sformatf("Buffer State: rd_ptr=%0d, pck_len_wr_ptr=%0d, pck_len_rd_ptr=%0d, empty=%0b, full=%0b, empty_de_assert=%0b, in_sop_r=%0b, in_sop_r1=%0b, in_sop_r2=%0b, in_eop_r=%0b, in_eop_r1=%0b, in_eop_r2=%0b",   
                 ref_rd_ptr, ref_pck_len_wr_ptr, ref_pck_len_rd_ptr, ref_buffer_empty, ref_buffer_full, ref_empty_de_assert, ref_in_sop_r, ref_in_sop_r1, ref_in_sop_r2, ref_in_eop_r, ref_in_eop_r1, ref_in_eop_r2), UVM_LOW)
        
        // No longer need buffer_empty_r since we use simple wr_lvl-based logic
        
        // Packet length buffer conditions
        ref_pck_len_full = (ref_pck_len_wr_ptr == ref_pck_len_rd_ptr) ? 0 :
                          (({~ref_pck_len_wr_ptr[5], ref_pck_len_wr_ptr[4:0]} == ref_pck_len_rd_ptr) ? 1 : 0);
        ref_pck_len_empty = (ref_pck_len_wr_ptr == ref_pck_len_rd_ptr) ? 1 : 0;
    endfunction
    
    function void update_write_level_next();
        // CRITICAL FIX: Write level is now calculated from pointers (wr_ptr - rd_ptr)
        // This function is kept for compatibility but wr_lvl_next is calculated in the final phase
        // RTL: wr_lvl = wr_ptr - rd_ptr
        
        if (ref_reset_active) begin
            // Hardware or software reset active: keep wr_lvl_next at 0 (matching RTL reset behavior)
            ref_wr_lvl_next = 0;
            `uvm_info("WR_LVL_DEBUG", $sformatf("Time=%0t: RESET ACTIVE: ref_wr_lvl_next kept at 0 (matching DUT reset behavior)", $time), UVM_LOW)
        end else begin
            // CRITICAL FIX: wr_lvl_next is calculated from pointers in the final phase
            // This ensures correct calculation: wr_lvl = wr_ptr - rd_ptr
            ref_wr_lvl_next = ref_wr_lvl;  // Keep current value, will be updated in final phase
        end
        
        // Debug wr_lvl calculation details
        `uvm_info("WR_LVL_DEBUG", $sformatf("wr_lvl_next placeholder: wr_en=%0b, rd_en=%0b, buffer_full=%0b, buffer_empty=%0b, current_wr_lvl=%0d, wr_ptr=%0d, rd_ptr=%0d", 
                 ref_wr_en, ref_rd_en, ref_buffer_full, ref_buffer_empty, ref_wr_lvl, ref_wr_ptr, ref_rd_ptr), UVM_LOW)
    endfunction

    function void update_internal_overflow();
        // Internal overflow logic (matching int_buffer_top's always_ff)
        // Use previous cycle's buffer states for calculation
        if (ref_buffer_full && ref_wr_en) begin
            ref_overflow = 1;
        end else begin
            ref_overflow = 0;
        end
    endfunction

    function void update_overflow_underflow(pkt_proc_seq_item tr);
        // CRITICAL FIX: Overflow detection should be delayed by 2 cycles to match DUT's registered output
        // DUT's pck_proc_overflow goes high AFTER one clock pulse after pck_proc_full goes high
        // Scoreboard should use two-cycle delayed buffer_full state to match DUT timing
        
        // Overflow detection - use two-cycle delayed buffer_full state
        if (tr.enq_req && ref_buffer_full_prev2) begin
            ref_pck_proc_overflow = 1;
            `uvm_info("OVERFLOW_DEBUG", $sformatf("Time=%0t: Overflow detected (delayed by 2 cycles): enq_req=%0b, buffer_full_prev2=%0b", 
                     $time, tr.enq_req, ref_buffer_full_prev2), UVM_LOW)
        end else begin
            ref_pck_proc_overflow = 0;
        end

        // Underflow detection - use previous cycle's buffer_empty state
        if (tr.deq_req && ref_buffer_empty_prev) begin
            ref_pck_proc_underflow = 1;
            `uvm_info("UNDERFLOW_DEBUG", $sformatf("Time=%0t: Underflow detected (delayed by 1 cycle): deq_req=%0b, buffer_empty_prev=%0b", 
                     $time, tr.deq_req, ref_buffer_empty_prev), UVM_LOW)
        end else begin
            ref_pck_proc_underflow = 0;
        end
        
    endfunction

    function void update_outputs(pkt_proc_seq_item tr);
        // Generate expected outputs
        ref_out_sop = 0;
        ref_out_eop = 0;
        
        // CRITICAL FIX: Scoreboard mirrors RTL exactly using present_state and deq_req_r
        // RTL uses present_state_r (current state after always_ff update) for output generation
        // Scoreboard must use the state that was active BEFORE the current cycle's state advance
        unique case (read_state_prev)  // ← Use previous state (matching RTL present_state_r timing)
            IDLE_R: begin
                ref_out_sop = 0;
                ref_out_eop = 0;
            end
            READ_HEADER: begin
                if (ref_deq_req_r) begin  // ← Use registered version (matching RTL)
                    ref_out_sop = 1;
                    ref_out_eop = 0;
                    // CRITICAL FIX: Don't increment count_r here - RTL does it in always_ff (next cycle)
                    // The output generation should use the current count_r value, not the incremented one
                    `uvm_info("COUNT_DEBUG", $sformatf("Time=%0t: READ_HEADER: out_sop=1, count_r=%0d (will increment to %0d next cycle)", 
                             $time, ref_count_r, ref_count_r + 1), UVM_LOW)
                end
            end
            READ_DATA: begin
                if (ref_deq_req_r) begin  // ← Use registered version (matching RTL)
                    // CRITICAL FIX: Check if this is the last beat BEFORE incrementing count_r
                    // This ensures out_eop is generated on the correct beat
                    if (ref_count_r == (ref_packet_length - 1)) begin
                        ref_out_eop = 1;
                        ref_count_r = 0; // packet boundary
                        `uvm_info("COUNT_DEBUG", $sformatf("Time=%0t: READ_DATA count_r reset to 0 (packet complete, length=%0d, was at %0d)", 
                                 $time, ref_packet_length, ref_count_r), UVM_LOW)
                    end else begin
                        ref_out_eop = 0;
                        // CRITICAL FIX: count_r increment is now handled in final updates (matching RTL always_ff)
                        `uvm_info("COUNT_DEBUG", $sformatf("Time=%0t: READ_DATA: out_eop=0, count_r=%0d (will increment to %0d next cycle)", 
                                 $time, ref_count_r, ref_count_r + 1), UVM_LOW)
                    end
                end
            end
        endcase
        
        // // Combinational output signals (matching RTL exactly)
        update_combinational_outputs(tr);
        
        // Debug out_sop calculation (now using previous state to match RTL timing)
        `uvm_info("OUT_SOP_DEBUG", $sformatf("out_sop/eop: prev_state=%0d, curr_state=%0d, deq_req_r=%0b, count_r=%0d, pck_len=%0d, out_sop=%0b, out_eop=%0b (using prev_state)", 
                 read_state_prev, read_state, ref_deq_req_r, ref_count_r, ref_packet_length, ref_out_sop, ref_out_eop), UVM_LOW)
        
        // Debug count_r timing alignment with RTL
        `uvm_info("COUNT_R_TIMING", $sformatf("Time=%0t: count_r timing: current=%0d, will_update=%0b, out_eop=%0b (RTL always_ff timing)", 
                 $time, ref_count_r, ref_deq_req_r && (read_state_prev == READ_HEADER || read_state_prev == READ_DATA), ref_out_eop), UVM_LOW)
        
        // Debug count_r priority logic to match RTL
        if (ref_out_eop) begin
            `uvm_info("COUNT_R_PRIORITY", $sformatf("Time=%0t: count_r PRIORITY: out_eop=1 takes precedence, count_r will be reset to 0", $time), UVM_LOW)
        end else if (ref_deq_req_r && (read_state_prev == READ_HEADER || read_state_prev == READ_DATA)) begin
            `uvm_info("COUNT_R_PRIORITY", $sformatf("Time=%0t: count_r PRIORITY: out_eop=0, count_r will increment from %0d to %0d", 
                     $time, ref_count_r, ref_count_r + 1), UVM_LOW)
        end
    endfunction

    function void update_combinational_outputs(pkt_proc_seq_item tr);
        // CRITICAL FIX: pck_proc_full should be based on wr_lvl, not pointer comparison
        // DUT logic: pck_proc_full = 1 when wr_lvl == DEPTH (buffer is full)
        // This matches the actual RTL behavior, not the complex pointer-based logic
        ref_buffer_full = (ref_wr_lvl == DEPTH) ? 1 : 0;  // Use parameter instead of hardcoded value
        
        // CRITICAL FIX: pck_proc_empty should be based on wr_lvl, not pointer comparison
        // DUT logic: pck_proc_empty = 1 when wr_lvl > 0 (buffer has data)
        // This matches the actual RTL behavior, not the complex pointer-based logic
        ref_buffer_empty = (ref_wr_lvl > 0) ? 0 : 1;
        
        // CRITICAL FIX: pck_proc_almost_full threshold should be DEPTH - almost_full_value
        // DUT logic: pck_proc_almost_full = 1 when wr_lvl >= (DEPTH - almost_full_value)
        // This matches the actual RTL behavior
        ref_pck_proc_almost_full = (ref_wr_lvl >= (DEPTH - tr.pck_proc_almost_full_value));
        
        // pck_proc_almost_empty (from buffer_almost_empty) - matching RTL assign
        // Use transaction value, not hardcoded value
        ref_pck_proc_almost_empty = (ref_wr_lvl <= tr.pck_proc_almost_empty_value);

    endfunction

    function void compare_outputs(pkt_proc_seq_item tr);
        // Debug information
        `uvm_info("SCOREBOARD_DEBUG", $sformatf("Time=%0d: DUT wr_lvl=%0d, ref_wr_lvl=%0d, DUT_empty=%0b, ref_empty=%0b, DUT_rd_data=0x%0h, ref_rd_data=0x%0h", 
                 $time, tr.pck_proc_wr_lvl, ref_wr_lvl, tr.pck_proc_empty, ref_buffer_empty, tr.rd_data_o, ref_rd_data_o), UVM_LOW)
        
        // Compare all outputs with reference model
        if (tr.out_sop !== ref_out_sop) begin
            `uvm_error("SCOREBOARD_NEW", $sformatf("out_sop mismatch: expected=%0b, got=%0b", ref_out_sop, tr.out_sop))
            errors++;
        end
        
        if (tr.out_eop !== ref_out_eop) begin
            `uvm_error("SCOREBOARD_NEW", $sformatf("out_eop mismatch: expected=%0b, got=%0b", ref_out_eop, tr.out_eop))
            errors++;
        end
        
        // CRITICAL FIX: Compare rd_data_o only when ref_deq_req_r is high (matching RTL timing)
        // RTL generates rd_data_o based on deq_req_r, not the current cycle's deq_req
        // CRITICAL FIX: Handle concurrent read/write operations properly
        bit data_available_for_comparison = 0;
        if (!ref_buffer_empty) begin
            // Normal case: data available in buffer
            data_available_for_comparison = 1;
        end else if (ref_wr_en && (ref_wr_ptr == ref_rd_ptr)) begin
            // Special case: writing to current read location, data will be available after write
            data_available_for_comparison = 1;
        end
        
        if (ref_deq_req_r && data_available_for_comparison) begin
            if (tr.rd_data_o !== ref_rd_data_o) begin
                `uvm_error("SCOREBOARD_NEW", $sformatf("rd_data_o mismatch: expected=0x%0h, got=0x%0h (deq_req_r=%0b, state=%0d)", 
                         ref_rd_data_o, tr.rd_data_o, ref_deq_req_r, read_state))
                errors++;
            end
        end
        
        if (tr.pck_proc_full !== ref_buffer_full) begin
            `uvm_error("SCOREBOARD_NEW", $sformatf("pck_proc_full mismatch: expected=%0b, got=%0b", ref_buffer_full, tr.pck_proc_full))
            errors++;
        end
        
        if (tr.pck_proc_empty !== ref_buffer_empty) begin
            `uvm_error("SCOREBOARD_NEW", $sformatf("pck_proc_empty mismatch: expected=%0b, got=%0b", ref_buffer_empty, tr.pck_proc_empty))
            errors++;
        end
        
        if (tr.pck_proc_almost_full !== ref_pck_proc_almost_full) begin
            `uvm_error("SCOREBOARD_NEW", $sformatf("pck_proc_almost_full mismatch: expected=%0b, got=%0b", ref_pck_proc_almost_full, tr.pck_proc_almost_full))
            errors++;
        end
        
        if (tr.pck_proc_almost_empty !== ref_pck_proc_almost_empty) begin
            `uvm_error("SCOREBOARD_NEW", $sformatf("pck_proc_almost_empty mismatch: expected=%0b, got=%0b", ref_pck_proc_almost_empty, tr.pck_proc_almost_empty))
            errors++;
        end
        
        if (tr.pck_proc_overflow !== ref_pck_proc_overflow) begin
            `uvm_error("SCOREBOARD_NEW", $sformatf("pck_proc_overflow mismatch: expected=%0b, got=%0b", ref_pck_proc_overflow, tr.pck_proc_overflow))
            errors++;
        end
        
        if (tr.pck_proc_underflow !== ref_pck_proc_underflow) begin
            `uvm_error("SCOREBOARD_NEW", $sformatf("pck_proc_underflow mismatch: expected=%0b, got=%0b", ref_pck_proc_underflow, tr.pck_proc_underflow))
            errors++;
        end
        
        if (tr.packet_drop !== ref_packet_drop) begin
            `uvm_error("SCOREBOARD_NEW", $sformatf("packet_drop mismatch: expected=%0b, got=%0b", ref_packet_drop, tr.packet_drop))
            errors++;
        end
        
        // if (tr.pck_proc_wr_lvl !== ref_wr_lvl) begin
        //     `uvm_error("SCOREBOARD_NEW", $sformatf("pck_proc_wr_lvl mismatch: expected=%0d, got=%0d (wr_en=%0b, rd_en=%0b, buffer_full=%0b, buffer_empty=%0b, overflow=%0b)", ref_wr_lvl, tr.pck_proc_wr_lvl, ref_wr_en, ref_rd_en, ref_buffer_full, ref_buffer_empty, ref_overflow))
        //     errors++;
        // end
    endfunction

    function void report_phase(uvm_phase phase);
        super.report_phase(phase);
        `uvm_info("SCOREBOARD_NEW", $sformatf("New Scoreboard Report: Total=%0d, Errors=%0d", total_transactions, errors), UVM_LOW)
    endfunction

endclass 
